library verilog;
use verilog.vl_types.all;
entity CodecConfig_vlg_vec_tst is
end CodecConfig_vlg_vec_tst;
