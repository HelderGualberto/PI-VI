--Codec system configuration i2c

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CodecConfig is 
	port(
		
	);
end CodecConfig;

ARCHITECTURE archconfig of CodecConfig is
	begin
	
end archconfig;