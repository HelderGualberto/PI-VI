library verilog;
use verilog.vl_types.all;
entity CODECSystem_vlg_vec_tst is
end CODECSystem_vlg_vec_tst;
