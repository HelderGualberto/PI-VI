library verilog;
use verilog.vl_types.all;
entity FFTDivider32_vlg_vec_tst is
end FFTDivider32_vlg_vec_tst;
