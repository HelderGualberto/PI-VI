library verilog;
use verilog.vl_types.all;
entity CodecConfig_vlg_sample_tst is
    port(
        SCLK            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end CodecConfig_vlg_sample_tst;
