library verilog;
use verilog.vl_types.all;
entity FFTDivider32_vlg_check_tst is
    port(
        CLKout          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FFTDivider32_vlg_check_tst;
