-- Sistema digital analogico
LIBRARY ieee;
USE ieee.std_logic_1164.all;

Entity DASystem IS
	port(
		DACDAT : IN BIT;
		DACCLK : IN BIT
	);
	
END DASystem;

ARCHITECTURE DAArch of DASystem is
	begin
end DAArch;
