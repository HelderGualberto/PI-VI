library verilog;
use verilog.vl_types.all;
entity CODECSystem_vlg_sample_tst is
    port(
        CPUCLK          : in     vl_logic;
        DAdata          : in     vl_logic_vector(15 downto 0);
        sampler_tx      : out    vl_logic
    );
end CODECSystem_vlg_sample_tst;
